`include "fetch.v"
`include "decode.v"


module processor()

endmodule